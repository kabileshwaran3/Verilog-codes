//Write a testbench for a blocking-assigned flip-flop—verify its output.
module ff_blocking(
    input clk,
    input rst,
    input d,
    output reg q);
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            q = 0;        
        end else begin
            q = d;
        end
    end
endmodule
