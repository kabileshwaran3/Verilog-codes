`timescale 1ns / 1ps

module implicit_or(input a,input b,   
                     output out);

    assign out=a|b;
endmodule
